*AXA3

.subckt AXA3 a b cin sum cout vdd
*DUT
    *PMOS
        Mp1 vdd a tmp vdd pmos_rvt nfin=n
        Mp2 tmp b xo vdd pmos_rvt nfin=n
        Mp3 gnd xo sum vdd pmos_rvt nfin=n
        Mp4 cin xo cout vdd pmos_rvt nfin=n
    *NMOS
        Mn1 xo b a gnd nmos_rvt nfin=n
        Mn2 xo a b gnd nmos_rvt nfin=n
        Mn3 cin xo sum gnd nmos_rvt nfin=n
        Mn4 a xo cout gnd nmos_rvt nfin=n
.ends
