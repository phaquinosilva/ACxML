* 8 bit comparator using subtractors

.include 8bRCA.cir

** A - B --- result of a > b in s7
.subckt 8b_sub_comp a0 a1 a2 a3 a4 a5 a6 a7 b0 b1 b2 b3 b4 b5 b6 b7 gt vdd
*********************************
**DUT
*inverters
Xb0 b0 nb0 vdd Inv
Xb1 b1 nb1 vdd Inv
Xb2 b2 nb2 vdd Inv
Xb3 b3 nb3 vdd Inv
Xb4 b4 nb4 vdd Inv
Xb5 b5 nb5 vdd Inv
Xb6 b6 nb6 vdd Inv
Xb7 b7 nb7 vdd Inv
*adders
Xadd a0 a1 a2 a3 a4 a5 a6 a7 nb0 nb1 nb2 nb3 nb4 nb5 nb6 nb7 vdd s0 s1 s2 s3 s4 s5 s6 gt vdd 8bRCA
********************************
.ends