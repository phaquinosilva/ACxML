** 4 bit binary reduced logic comparator

* XNOR
.subckt xnor a b out vdd
Mpa vdd a ab a pmos_rvt nfin=3
Mpb ab b out b pmos_rvt nfin=3
Mna out a b a nmos_rvt nfin=3
Mnb out b a b nmos_rvt nfin=3
.ends

.subckt nand2 a b out vdd
Mpa vdd a out a pmos_rvt nfin=3
Mpb vdd b out b pmos_rvt nfin=3
Mna out a ab a nmos_rvt nfin=3
Mnb ab b gnd b nmos_rvt nfin=3
.ends

.subckt nand3 a b c out vdd
Mpa vdd a out a pmos_rvt nfin=3
Mpb vdd b out b pmos_rvt nfin=3
Mpc vdd c out c pmos_rvt nfin=3
Mna out a ab a nmos_rvt nfin=3
Mnb ab b bc b nmos_rvt nfin=3
Mnb bc c gnd c nmos_rvt nfin=3
.ends

.subckt nor2 a b out vdd
Mpa vdd a ab a pmos_rvt nfin=3
Mpb ab b out b pmos_rvt nfin=3
Mna out a gnd a nmos_rvt nfin=3
Mnb out b gnd b nmos_rvt nfin=3
.ends

.subckt nand4 a b c d out vdd
Xn20 a b n0 vdd nand2
Xn21 c d n1 vdd nand2
Xo n0 n1 nout vdd nor2
Xinv nout out vdd Inv
.ends

.subckt nand5 a b c d e out vdd
Xn2 a b n0 vdd nand2
Xn3 c d e n1 vdd nand3
Xo n0 n1 nout vdd nor2
Xinv nout out vdd Inv
.ends

* result of a > b in s3
.subckt 4b_ded_comp a0 a1 a2 a3 b0 b1 b2 b3 geq vdd
*DUT
* A xnor B
Xeq1 a1 b1 eq1 vdd xnor
Xeq2 a2 b2 eq2 vdd xnor
Xeq3 a3 b3 eq3 vdd xnor

* not A
Xa0 a0 na0 vdd Inv
Xa1 a1 na1 vdd Inv
Xa2 a2 na2 vdd Inv
Xa3 a3 na3 vdd Inv

* greater
Xn3 b3 na3 n3 vdd nand2
Xn2 b2 na2 eq3 n2 vdd nand3
Xn1 b1 na1 eq3 eq2 n1 vdd nand4
Xn0 b0 na0 eq3 eq2 eq1 n0 vdd nand5

Xgeq n3 n2 n1 n0 geq vdd nand4

.ends