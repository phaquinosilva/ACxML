**inverter

*circuit - inverter
.subckt inv in out vdd
  Mp vdd in out in pmos_rvt nfin=n
  Mn out in gnd in nmos_rvt nfin=n
.ends
