*AMA2 validation

*model
.include 7nm_FF.pm

*param
.param vdd = 0.7V
.param n = 3
.option post = 2

*sources
Vvdut vdut gnd vdd
Vvdd1 vdd1 gnd vdd
* Vvdd2 vdd2 gnd vdd
*validation sources
Va a_in gnd PWL(0n vdd)
Vb b_in gnd PWL(0n 0)
Vcin c_in gnd PWL(0n vdd)

.include inverter.cir
.include fas/ama2.cir

*IN fanout
Xinv1 a_in a_in1 vdd1 Inv
Xinv2 a_in1 a vdd1 Inv

Xinv3 b_in b_in1 vdd1 Inv
Xinv4 b_in1 b vdd1 Inv

Xinv5 c_in c_in1 vdd1 Inv
Xinv6 c_in1 cin vdd1 Inv

*****************DUT******************
XDUT a b cin sum cout vdut AMA2

*OUT fanout
Csum sum gnd 1f
Ccout cout gnd 1f

*simulation
.tran 0.1ns 2ns

.end

