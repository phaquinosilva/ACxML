
* predition model
.include 7nm_FF.cir

* technology specific
.param vdd = 0.7V
.param n = 3

* output formatting - cscope and csv
.option post = 2
.option measform = 3

* default voltage sources used
Vvdd1 vdd1 gnd vdd
Vvdut vdut gnd vdd
* Vvdd2 vdd2 gnd vdd

