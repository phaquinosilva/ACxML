**inverter

*circuit - inverter
.subckt Inv in out vdd
  Mp vdd in out in pmos_rvt nfin=3
  Mn out in gnd in nmos_rvt nfin=3
.ends
