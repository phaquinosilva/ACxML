*** MODELO ***

**modelo preditivo
.include __.pm

.include param.cir

** fontes
Vvdut vdut gnd vdd
Vvdd1 vdd1 gnd vdd
Vvdd2 vdd2 gnd vdd

*incluir arquivo de entradas
.include sources.cir

** incluir modelo de somador
.include ..

**descricao circuito
*load
..
*DUT
..
*FO4
..

** measures
*energia
.measure carga load
.measure carga DUT
.measure carga FO4
*atraso
.measure todos os atrasos
..

** tipo de simulação
.tran ..

.end
