**MIRROR

.subckt EMA a b cin sum cout vdd
*DUT
    *PMOS
        Mp1 vdd a t1 a pmos_rvt l=len nfin=n
        Mp2 vdd b t1 b pmos_rvt l=len nfin=n
        Mp3 t1 cin co cin pmos_rvt l=len nfin=n
        Mp4 vdd b ta b pmos_rvt l=len nfin=n
        Mp5 ta a co a pmos_rvt l=len nfin=n
        Mp6 vdd a t2 a pmos_rvt l=len nfin=n
        Mp7 vdd b t2 b pmos_rvt l=len nfin=n
        Mp8 vdd cin t2 cin pmos_rvt l=len nfin=n
        Mp9 t2 co su co pmos_rvt l=len nfin=n
        Mpa vdd a tb a pmos_rvt l=len nfin=n
        Mpb tb b tc b pmos_rvt l=len nfin=n
        Mpc tc cin su cin pmos_rvt l=len nfin=n
    *NMOS
        Mn1 co cin t3 cin nmos_rvt l=len nfin=n
        Mn2 t3 a gnd a nmos_rvt l=len nfin=n
        Mn3 t3 b gnd b nmos_rvt l=len nfin=n
        Mn4 co a tb1 a nmos_rvt l=len nfin=n
        Mn5 tb1 b gnd b nmos_rvt l=len nfin=n
        Mn6 su co t4 co nmos_rvt l=len nfin=n
        Mn7 t4 a gnd a nmos_rvt l=len nfin=n
        Mn8 t4 b gnd b nmos_rvt l=len nfin=n
        Mn9 t4 cin gnd cin nmos_rvt l=len nfin=n
        Mnb tb2 b ta2 b nmos_rvt l=len nfin=n
        Mna su cin tb2 cin nmos_rvt l=len nfin=n
        Mnc ta2 a gnd a nmos_rvt l=len nfin=n

    *inverters for accurate results
        Xsum su sum vdd gnd Inv
        Xcout co cout vdd gnd Inv
.ends
