*AMA1

.subckt AMA1 a b cin sum cout vdd
*DUT
    *PMOS
        Mp1 vdd b sc1 b pmos_rvt nfin=n
        Mp2 sc1 cin co cin pmos_rvt nfin=n
        Mp3 vdd b sc2 b pmos_rvt nfin=n
        Mp4 sc2 a co a pmos_rvt nfin=n
        Mp5 vdd co tmp1 co pmos_rvt nfin=n
        Mp6 vdd tmp1 sum tmp1 pmos_rvt nfin=n
    *NMOS
        Mn1 co cin sd1 cin nmos_rvt nfin=n
        Mn2 sd1 a gnd a nmos_rvt nfin=n
        Mn3 co b gnd b nmos_rvt nfin=n
        Mn4 tmp1 co gnd co nmos_rvt nfin=n
        Mn5 sum tmp1 gnd tmp1 nmos_rvt nfin=n
    *inverter for correct output
        Xcout co cout vdd Inv
.ends
