**inverter

*circuit - inverter
.subckt Inv in out vdd
  Mp vdd in out in pmos_rvt L=len nfin=n
  Mn out in gnd in nmos_rvt L=len nfin=n
.ends
