*** MODELO ***

**modelo preditivo
.include ..

** parametros (predefinidos para FinFET)
.param vdd = 0.7V
.param len = 7nm
*numero de fins
.param n = 3
.option post = 2
*define saída em .csv
.option measform= 3

** fontes
Vvdut vdut gnd vdd
Vvdd1 vdd1 gnd vdd
Vvdd2 vdd2 gnd vdd
*incluir arquivo de entradas
.include ..

** incluir modelo de somador
.include ..

**descricao circuito
*load
..
*DUT
..
*FO4
..

** measures
*energia
.measure carga load
.measure carga DUT
.measure carga FO4
*atraso
.measure todos os atrasos
..

** tipo de simulação
.tran ..

.end
